`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2025/05/02 13:32:28
// Design Name: 
// Module Name: wechat_jump_fsm
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////
module wechat_jump_fsm (
    // ???????????
    input  wire        clk_machine,    // ????? (25.175MHz)
    input  wire        rst_machine,    // ????�� (????��)
    input  wire        i_btn,          // ??????????
    input  wire        i_btn_origin,

    //??jump????????
    input  wire        i_jump_done,    // ?????????????????
    input  wire [10:0] i_jump_dist,
    input  wire [8:0] i_jump_height,
    output wire  [10:0]  o_jump_v_init,  // ????????
    output reg         o_jump_en,       // ???????????
    
    
    // ?????
    output reg  [2:0]  state,          // ???????
    
    // ????????graphics???????
    output reg  [10:0] o_x_man,
    output reg  [10:0] o_y_man,
    output reg  [10:0] o_x_block1,     // ????1??X????
    output reg  [10:0] o_x_block2,     // ????2??X????
    output reg         o_en_block2,     // ????2??????
    output reg  [3:0]  o_type_block1, // ????1????
    output reg  [3:0]  o_type_block2, // ????2????
    //???????????????color?????type?????graphics??block?��???????????????????????
    //??????????????��??��??0~5
    output wire  [3:0]  o_squeeze_man,  // ��?????? (0-14)

    //??????????????graphics??�?????????????????????????
    output reg o_title,
    output reg o_gameover,

    output reg  [9:0] o_score,         // ?��?

    output reg o_perfect
    
    );

    // ================= ?????? ================= //
    localparam INIT = 3'd0;  // ??????? (????��?????)
    localparam RELD = 3'd1;  // ?????��????
    localparam WAIT = 3'd2;  // ?????????
    localparam ACCU = 3'd3;  // ??????
    localparam JUMP = 3'd4;  // ???????
    localparam LAND = 3'd5;  // ????��???
    localparam OVER = 3'd6;  // ?????????

    // ================= ???????? ================= //
    //????��??????
    localparam ORIGIN         = 32'd0;   // ??????????
    localparam ORIGIN_STARTUP = 32'd100;     // INIT?????????1?????????????
    localparam BLOCK_WIDTH    = 32'd35;   // ????????????????��??????????????��????????��??????????
    localparam BLOCK_CENTER_WIDTH = 32'd10; // ???????????
    localparam BLOCK2_OFFSET  = 32'd180;    // ????2?????????
    localparam MAX_SQUEEZE    = 4'd14;     // ???????????????????��??0-14

    // ================= ?????? ================= //
    reg  [16:0] cnt_clk_reload;       // ??��??????????
    reg  [31:0] cnt_v_init;           // ????????????????cnt_v_init???????????????clk??????
    /*????????��???????????��?????????��????????????????????????????????????��??????*/
    reg         reload_done;          // ??��?????
    wire [6:0]  random;               // ???????random?????????????
    reg new_game;                     // ?????��?????????????????????????????????

    reg  [10:0] relative_x;           // ??????????????��???????


    // ??????
    assign o_jump_v_init = cnt_v_init[24:18];  // ?cnt_v_init?????7��???????????��??0-127??jump????��?????127??????????256???????260
    assign o_squeeze_man = state==JUMP? 0 : cnt_v_init[24:18]*14/127%15;   // ?cnt_v_init?????4��??????????��??0-14?????????15???��???????



    // ================= ???????? ================= //
    //??????????????��?
    always @(posedge clk_machine or posedge rst_machine) begin
        if (rst_machine) begin           // ??��?????��?
            state <= RELD;               // ????��??????
            new_game       <= 1'b1;     //rst_machine???????????????????
            o_title        <= 1'b1; 
            o_gameover     <= 1'b0;
            o_jump_en      <= 1'b0;
            o_score        <= 10'd0;
            
            relative_x <= 11'd0;                 // ???????????
            o_perfect     <= 1'b0;
        end else begin                 // ??��???????
            case (state)
                INIT: begin              
                    state <= RELD;           // INIT????????RELD??
                end
                RELD: begin             // RELD?????????1????????��??
                    if(new_game) begin  // ???????????????????????????
                        o_title <= 1'b1;
                    end
                    if (reload_done || o_x_block1==ORIGIN) begin // ??��???????????????��??????
                        state <= WAIT;      // ????????????
                    end else begin
                        state <= RELD;      // ????��??��????????��????
                    end
                end
                WAIT: begin             // ?????????
                    if (i_btn) begin       // ?????��????????????????
                        state <= ACCU; 
                        if(new_game) begin
                            new_game <= 1'b0;   //??��??????????????????????
                            o_title <= 1'b0;   // ?????????
                        end
                    end
                end
                ACCU: begin             // ??????
                    if (i_btn) begin    //???��?????????????????????
                        state <= ACCU;
                    end else begin
                        o_jump_en=1'b1;
                        state <= JUMP;  //??????????????????
                    end
                end
                JUMP: begin             // ???????
                    if (i_jump_done) begin // ?????????????????????????��???
                        o_jump_en=1'b0;
                        state <= LAND;
                    end else begin
                        state <= JUMP;      // ???????????????????????
                    end
                end
                LAND: begin             // ????��???
                    if (o_x_man <= BLOCK_WIDTH) begin // ��??��?????????
                        state <= WAIT;      // ??????��??????
                    end else if((o_x_man < o_x_block2)?
                        (o_x_block2-o_x_man <BLOCK_CENTER_WIDTH)
                        :(o_x_man-o_x_block2 <BLOCK_CENTER_WIDTH)) begin
                        o_score <= o_score + 2; // ?��??2
                        o_perfect <= 1'b1;
                        relative_x <= 0;
                        state <= INIT;      // ????��?????
                    end else if((o_x_man < o_x_block2)?
                        (o_x_block2-o_x_man <BLOCK_WIDTH)
                        :(o_x_man-o_x_block2 <BLOCK_WIDTH)) begin
                        o_score <= o_score + 1; // ?��??1
                        o_perfect <= 1'b0;
                        relative_x <= o_x_man - o_x_block2; // ??????????????????��???????,????��??????????????????��?��???
                        state <= INIT;      // ????��?????
                    end else begin
                        state <= OVER;      // ?????????
                    end
                end
                OVER: begin             // ?????????
                    state <= OVER;          // ????????
                    o_gameover <= 1'b1;    // ??????????????
                end
                default: begin           // ??????
                    state <= RELD;          // ??????????
                end
            endcase
        end
    end

    /*????????��???????always????��?????????*/
    
    //????????????????
    random #(7) random_inst (
        .clk_random(clk_machine),
        .rst_random(rst_machine),
        .i_roll(i_btn_origin),
        .o_random_binary(random)
    );

    //????????????��???
    always @(posedge clk_machine or posedge rst_machine) begin
        if (rst_machine) begin
            o_x_block1 <= ORIGIN_STARTUP;     // ??????1??????2??????ORIGIN_STARTUP??��??
            o_x_block2 <= ORIGIN_STARTUP;     
            o_en_block2 <= 1'b0;              // ????????2
            reload_done <= 1'b0;             
            cnt_clk_reload <= 17'd0;          // ??��??????????
        end else begin
            case (state)
                INIT: begin
                    cnt_clk_reload <= 17'd0;
                    o_x_block1 <= o_x_block2;    // ????��?????
                    o_x_block2 <= o_x_block2;    // ????��?��???
                    o_en_block2 <= 1'b0;
                    reload_done <= 1'b0;
                end
                RELD: begin
                    if(o_x_block1 > ORIGIN) begin       // ??????1??????????ORIGIN��??
                        if (cnt_clk_reload == 17'h1ffff) begin // ?????clk_machine????13?��??
                            cnt_clk_reload <= 17'd0; // ??��??????
                            o_x_block1 <= o_x_block1 - 1; // ????????1
                        end else begin
                            cnt_clk_reload <= cnt_clk_reload + 1; // ????????1
                            o_x_block1 <= o_x_block1; // ????1��?��???
                        end
                        o_x_block2 <= o_x_block2;
                        o_en_block2 <= 1'b0;
                        reload_done <= 1'b0;
                    end else begin                    // ??????1????????ORIGIN��??
                        cnt_clk_reload <= 17'd0;
                        o_x_block1 <= ORIGIN; // ??��????1
                        o_x_block2 <= ORIGIN + random + BLOCK2_OFFSET; // ??????????????????????????2??��??????
                        o_en_block2 <= 1'b1; // ???????2
                        reload_done <= 1'b1; // ??��??????
                    end
                end
                default: begin
                    cnt_clk_reload <= 17'd0;
                    o_x_block1 <= o_x_block1;     // ???????
                    o_x_block2 <= o_x_block2;     // ???????
                    o_en_block2 <= o_en_block2;      // ?????????
                    reload_done <= 1'b0;             // ??��??????
                end
            endcase
        end
    end
    
    // ????????????��???
    always@(posedge clk_machine or posedge rst_machine) begin
        if(rst_machine) begin
            o_type_block1 <= 5'd5;
            o_type_block2 <= 5'd0;
        end else begin
            case(state) 
                INIT:begin
                    o_type_block1 <= o_type_block2;
                    if(o_type_block2 == 5) begin        //??????????��??0~5
                        o_type_block2 <= 0;
                    end else begin
                        o_type_block2 <= o_type_block2 + 1;
                    end 
                end 
                
                default:begin
                    o_type_block1 <= o_type_block1;
                    o_type_block2 <= o_type_block2;
                end 
            endcase
        end
    end
    
    //????????????��??????????
    always @(posedge clk_machine or posedge rst_machine) begin
        if (rst_machine) begin
            cnt_v_init <= 0;
        end else begin
            case(state)
                ACCU: begin
                    if (i_btn && cnt_v_init < 25'h1ffffff) begin //????cnt_v_init???????????????clk??????
                        cnt_v_init <= cnt_v_init + 1;
                    end else begin
                        cnt_v_init <= cnt_v_init;
                    end
                end
                JUMP: begin
                    if (i_jump_done) begin
                        cnt_v_init <= 0;
                    end else begin
                        cnt_v_init <= cnt_v_init;
                    end
                end
            endcase
        end
    end

    // ???��?????
    always@(posedge clk_machine or posedge rst_machine) begin
        if(rst_machine) begin
            o_x_man <= ORIGIN_STARTUP;
            o_y_man <= 0;
        end else begin
            case (state)
                INIT: begin
                    o_x_man <= o_x_man;
                    o_y_man <= 0;
                end

                RELD: begin
                    o_x_man <= o_x_block1 + relative_x;
                    o_y_man <= 0;
                end
                
                ACCU: begin
                    o_x_man <= o_x_man;
                    o_y_man <= 0;
                end
                
                JUMP: begin
                    o_x_man <= o_x_block1 + relative_x + i_jump_dist*400/260; //?????????????400     
                    o_y_man <= i_jump_height;       
                end
                
                LAND, OVER: begin
                    o_x_man <= o_x_man;
                    o_y_man <= 0;
                end
                

            endcase
        end
    end
            
    


endmodule