/******************************************************************************
 ** Logisim-evolution goes FPGA automatic generated Verilog code             **
 ** https://github.com/logisim-evolution/                                    **
 **                                                                          **
 ** Component : clkdiv                                                       **
 **                                                                          **
 *****************************************************************************/

module clkdiv( clk,
               div_res,
               rst );

   /*******************************************************************************
   ** The inputs are defined here                                                **
   *******************************************************************************/
   input clk;
   input rst;

   /*******************************************************************************
   ** The outputs are defined here                                               **
   *******************************************************************************/
   output reg [31:0] div_res;

   /*******************************************************************************
   ** The module functionality is described here                                 **
   *******************************************************************************/

   /*******************************************************************************
   ** Here all output connections are defined                                    **
   *******************************************************************************/
 always @(posedge clk) begin
     if(rst==1'b1) begin
         div_res<=32'b0;
     end
     else begin
         div_res<=div_res+32'b1;
     end
   end
endmodule
